// Quantization_tb.v

module Quantization_tb();

Quantization #(
  .INPUT_INTEGER_WIDTH(),
  .INPUT_DECIMAL_WIDTH(),
  .OUTPUT_INTEGER_WIDTH(),
  .OUTPUT_DECIMAL_WIDTH()
)


endmodule;